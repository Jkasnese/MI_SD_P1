
module nios_project (
	btn_external_connection_export,
	clk_clk,
	leds_external_connection_export);	

	input		btn_external_connection_export;
	input		clk_clk;
	output	[3:0]	leds_external_connection_export;
endmodule
